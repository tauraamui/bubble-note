module main

const emoji_pallette = [
	"⚠️", "🚨", "✨", "✅", "⭐"
]


// have season specific emojis
// const season_emoji_pallette = ["🎄"]


