module main

const emoji_pallette = [
	"⚠️", "🚨", "U+1f47e", "U+1f4a5", "U+1f624"
]


